library verilog;
use verilog.vl_types.all;
entity fpu_tb is
    generic(
        FLOAT_2_759     : integer := 1076919009;
        FLOAT_NEG3_875  : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        FLOAT_0_000663  : integer := 976098427;
        FLOAT_10_2283   : integer := 1092854743;
        OP_ADD          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        OP_SUB          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        OP_MUL          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        OP_DIV          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        OP_MIN          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        OP_MAX          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        OP_SQRT         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        OP_FEQ          : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        OP_FLT          : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        OP_FLE          : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        OP_CVT_WS       : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        OP_CVT_WUS      : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi1);
        OP_CVT_SW       : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        OP_CVT_SWU      : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of FLOAT_2_759 : constant is 1;
    attribute mti_svvh_generic_type of FLOAT_NEG3_875 : constant is 1;
    attribute mti_svvh_generic_type of FLOAT_0_000663 : constant is 1;
    attribute mti_svvh_generic_type of FLOAT_10_2283 : constant is 1;
    attribute mti_svvh_generic_type of OP_ADD : constant is 1;
    attribute mti_svvh_generic_type of OP_SUB : constant is 1;
    attribute mti_svvh_generic_type of OP_MUL : constant is 1;
    attribute mti_svvh_generic_type of OP_DIV : constant is 1;
    attribute mti_svvh_generic_type of OP_MIN : constant is 1;
    attribute mti_svvh_generic_type of OP_MAX : constant is 1;
    attribute mti_svvh_generic_type of OP_SQRT : constant is 1;
    attribute mti_svvh_generic_type of OP_FEQ : constant is 1;
    attribute mti_svvh_generic_type of OP_FLT : constant is 1;
    attribute mti_svvh_generic_type of OP_FLE : constant is 1;
    attribute mti_svvh_generic_type of OP_CVT_WS : constant is 1;
    attribute mti_svvh_generic_type of OP_CVT_WUS : constant is 1;
    attribute mti_svvh_generic_type of OP_CVT_SW : constant is 1;
    attribute mti_svvh_generic_type of OP_CVT_SWU : constant is 1;
end fpu_tb;
